module restador4bits ( 
	a,
	b,
	borrowin,
	difference,
	borrowout
	) ;

input [3:0] a;
input [3:0] b;
input  borrowin;
inout [3:0] difference;
inout  borrowout;
