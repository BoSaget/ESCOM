module cto ( 
	a,
	b,
	c,
	d,
	validado
	) ;

input  a;
input  b;
input  c;
input  d;
inout  validado;
