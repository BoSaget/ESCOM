module reg4 ( 
	d,
	clk,
	en,
	q
	) ;

input [3:0] d;
input  clk;
input  en;
inout [3:0] q;
