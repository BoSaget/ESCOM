module led ( 
	switch,
	leds
	) ;

input [3:0] switch;
inout [9:0] leds;
