module contador0_7 ( 
	t,
	clk,
	q,
	nq
	) ;

input  t;
input  clk;
inout [2:0] q;
inout [2:0] nq;
