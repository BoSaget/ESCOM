module multiplexor4_1 ( 
	control,
	entradas,
	salida
	) ;

input [1:0] control;
input [3:0] entradas;
inout  salida;
