module decodificador ( 
	dato,
	segmento
	) ;

input [3:0] dato;
inout [6:0] segmento;
